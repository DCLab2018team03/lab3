
module AudioConfig (
	clk_clk,
	reset_reset_n,
	audio_and_video_config_0_external_interface_SDAT,
	audio_and_video_config_0_external_interface_SCLK);	

	input		clk_clk;
	input		reset_reset_n;
	inout		audio_and_video_config_0_external_interface_SDAT;
	output		audio_and_video_config_0_external_interface_SCLK;
endmodule
