
module AudioCoreInterpolation(
    input   [15:0]  i_data_prev,
    input   [15:0]  i_data,
    input   [3:0]   i_divisor,
    output  [15:0]  o_quotient
);
endmodule